module router_top(input clock,resetn,read_enb_0,read_enb_1,read_enb_2,input [7:0]data_in,input pkt_valid,output [7:0]data_out_0,data_out_1,data_out_2,
		output valid_out_0,valid_out_1,valid_out_2,error,busy);
		wire [2:0] write_enb;
		wire detect_add,write_enb_reg,full_0,full_1,full_2,empty_0,empty_1,empty_2,soft_reset_0,soft_reset_1,soft_reset_2;
		wire fifo_full,parity_done,low_pkt_valid,lfd_state,ld_state,laf_state,full_state,rst_int_reg;
		wire [7:0] data_out;


		router_sync dut1(detect_add,write_enb_reg,clock,resetn,read_enb_0,read_enb_1,read_enb_2,empty_0,empty_1,empty_2,
				full_0,full_1,full_2,data_in[1:0],soft_reset_0,soft_reset_1,soft_reset_2,fifo_full,write_enb,valid_out_0,	
				valid_out_1,valid_out_2);
		router_fsm  controller_dut(clock,resetn,pkt_valid,parity_done,soft_reset_0,soft_reset_1,soft_reset_2,fifo_full,low_pkt_valid,	
					empty_0,empty_1,empty_2,data_in[1:0],busy,lfd_state,detect_add,ld_state,laf_state,
					full_state,write_enb_reg,rst_int_reg);
		router_reg register_dut(clock,resetn,pkt_valid,data_in,fifo_full,rst_int_reg,detect_add,ld_state,laf_state,full_state,lfd_state,
					parity_done,low_pkt_valid,error,data_out);
		router_fifo fifo_0(clock,resetn,write_enb[0],soft_reset_0,read_enb_0,lfd_state,data_out,empty_0,full_0,data_out_0);
		router_fifo fifo_1(clock,resetn,write_enb[1],soft_reset_1,read_enb_1,lfd_state,data_out,empty_1,full_1,data_out_1);
		router_fifo fifo_2(clock,resetn,write_enb[2],soft_reset_2,read_enb_2,lfd_state,data_out,empty_2,full_2,data_out_2);
			
endmodule